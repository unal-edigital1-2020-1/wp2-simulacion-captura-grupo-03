`timescale 10ns / 1ns
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:14:22 12/02/2019 
// Design Name: 
// Module Name:    cam_read 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module cam_read #(
		parameter AW = 15,  // Cantidad de bits  de la direcci�n
		parameter DW = 12   //tamaño de la data 
		)
		(
		CAM_px_data,  //estrada de los datos de la camara
		CAM_pclk,     //reloj 
		CAM_vsync,    //Señal Vsync para captura de datos
		CAM_href,	// Señal Href para la captura de datos
		rst,		//reset
		
		DP_RAM_regW, 	//Control de esctritura
		DP_RAM_addr_in,	//Dirección de memoria de entrada
		DP_RAM_data_in	//Data de entrada a la RAM
   );
	
	input [7:0] CAM_px_data;	//Data RGB 444 de la camara
		input CAM_pclk;		//Reloj de la camara
		input CAM_vsync;	//señal vsync de la camara
		input CAM_href;		//señal href de la camara
		input rst;		//reset de la camara 
		
		output reg DP_RAM_regW; 		//Registro del control de escritura 
	output reg [AW-1:0] DP_RAM_addr_in;	// Registro de salida de la dirección de memoria de entrada 
	output reg [DW-1:0] DP_RAM_data_in;	// Registro de salida de la data a escribir en memoria


//Maquina de estados	
	
parameter INIT=0,BYTE1=1,BYTE2=2,NOTHING=3,imaSiz=19199;
reg [1:0]status=0;

always @(posedge CAM_pclk)begin
    if(rst)begin
    status<=0;
     DP_RAM_data_in<=0;
     DP_RAM_addr_in<=0;
     DP_RAM_regW<=0;
    end
    else begin
	    
     case (status)
         INIT:begin 
		 	if(~CAM_vsync&CAM_href)begin // Cuando la señal vsync es 0 y href 1, se empieza con la escritura de los datos en memoria.
                	status<=BYTE2;
			 		DP_RAM_data_in[11:8]<=CAM_px_data[3:0]; // Se asignan los 4 bits menos significativos de la información que da la camara a los 4 bits mas significativos del dato a escribir
            end
         	else begin
                	DP_RAM_data_in<=0;
                	DP_RAM_addr_in<=0;
                	DP_RAM_regW<=0; 
         	end 
        end
         
         BYTE1:begin
		 DP_RAM_regW<=0; 					//Desactiva la escritura en memoria 
		 if(CAM_href)begin					//si la señal Href esta arriva, evalua si ya llego a la ultima posicion en memoria
                	if(DP_RAM_addr_in==imaSiz) 	DP_RAM_addr_in<=0;			//Si ya llego al final, reinicia la posición en memoria. 
                	else DP_RAM_addr_in<=DP_RAM_addr_in+1;	//Si aun no ha llegado a la ultima posición sigue recorriendo los espacios en memoria y luego escribe en ellos cuan do pasa al estado Byte2
                DP_RAM_data_in[11:8]<=CAM_px_data[3:0];
                status<=BYTE2;
         end
         else status<=NOTHING;   
         end
         
         BYTE2:begin							//En este estado se habilita la escritura en memoria
             	DP_RAM_data_in[7:0]<=CAM_px_data;
             	DP_RAM_regW<=1;    
             	status<=BYTE1;
         end
         
         NOTHING:begin						// es un estado de trnsición 	
             
			if(CAM_href)begin					// verifica la señal href y se asigna los 4 bits mas significativos y se mueve una posición en memoria
					status<=BYTE2;
					DP_RAM_data_in[11:8]<=CAM_px_data[3:0];
					DP_RAM_addr_in<=DP_RAM_addr_in+1;
			end
			else if (CAM_vsync) status<=INIT;		// Si vsync esta arriba inicializa la maquina de estados   
         end
         
		 default: status<=INIT;
    endcase
 end
end
		

/********************************************************************************

Por favor colocar en este archivo el desarrollo realizado por el grupo para la 
captura de datos de la camara 

debe tener en cuenta el nombre de las entradas  y salidad propuestas 

********************************************************************************/

endmodule
